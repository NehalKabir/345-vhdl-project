-------------------------------------------------------------------------------
--
-- Title       : ese 345 project part 1
-- Design      : ese 345 project part 1
-- Author      : Nehal Kabir and Thomas Plourde
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : D:\ESE382\half_adder\half_adder\src\half_adder.vhd
-- Generated   : Wed Feb  9 09:44:48 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {half_adder} architecture {half_adder}}

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity reg_file is
	 port(
	  reg1 :in std_logic_vector (127 downto 0);  
	 reg2 :in std_logic_vector (127 downto 0);
	 reg3 :in std_logic_vector (127 downto 0);
	 reg4 :in std_logic_vector (127 downto 0);
	 reg5 :in std_logic_vector (127 downto 0);
	 reg6 :in std_logic_vector (127 downto 0);
	 reg7 :in std_logic_vector (127 downto 0);
	 reg8 :in std_logic_vector (127 downto 0);
	 reg9 :in std_logic_vector (127 downto 0);
	 reg10 :in std_logic_vector (127 downto 0);
	 reg11 :in std_logic_vector (127 downto 0);
	 reg12 :in std_logic_vector (127 downto 0);
	 reg13 :in std_logic_vector (127 downto 0);
	 reg14 :in std_logic_vector (127 downto 0);
	 reg15 :in std_logic_vector (127 downto 0);
	 reg16 :in std_logic_vector (127 downto 0);
	 reg17 :in std_logic_vector (127 downto 0);
	 reg18 :in std_logic_vector (127 downto 0);
	 reg19 :in std_logic_vector (127 downto 0);
	 reg20 :in std_logic_vector (127 downto 0);
	 reg21 :in std_logic_vector (127 downto 0);
	 reg22 :in std_logic_vector (127 downto 0);
	 reg23 :in std_logic_vector (127 downto 0);
	 reg24 :in std_logic_vector (127 downto 0);
	 reg25 :in std_logic_vector (127 downto 0);
	 reg26 :in std_logic_vector (127 downto 0);
	 reg27 :in std_logic_vector (127 downto 0);
	 reg28 :in std_logic_vector (127 downto 0);
	 reg29 :in std_logic_vector (127 downto 0);
	 reg30 :in std_logic_vector (127 downto 0);
	 reg31 :in std_logic_vector (127 downto 0);
	 reg32 :in std_logic_vector (127 downto 0);

	 write_reg :in std_logic_vector (127 downto 0);
	 
	 output1 : out std_logic_vector (127 downto 0);
	 output2 : out std_logic_vector (127 downto 0);
	 output3 : out std_logic_vector (127 downto 0)
	 
	     );
end reg_file;

--}} End of automatically maintained section

architecture reg_file of reg_file is
signal write: std_logic;
begin

	 -- enter your statements here --

end reg_file;
