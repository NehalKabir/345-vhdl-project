-------------------------------------------------------------------------------
--
-- Title       : instruction_buffer
-- Design      : project_part1
-- Author      : thomas plourde
-- Company     : HP Inc.
--
-------------------------------------------------------------------------------
--
-- File        : E:\ESE 345\Project_attempt2\project_part1\src\instruction_buffer.vhd
-- Generated   : Sun Nov 13 15:16:38 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {instruction_buffer} architecture {instruction_buffer}}

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity instruction_buffer is
port(
	r1 :in std_logic_vector (24 downto 0);	  
	r2 :in std_logic_vector (24 downto 0);
	r3 :in std_logic_vector (24 downto 0);
	r4 :in std_logic_vector (24 downto 0);
	r5 :in std_logic_vector (24 downto 0);
	r6 :in std_logic_vector (24 downto 0);
	r7 :in std_logic_vector (24 downto 0);
	r8 :in std_logic_vector (24 downto 0);
	r9 :in std_logic_vector (24 downto 0);
	r10 :in std_logic_vector (24 downto 0);	   
	
	r11 :in std_logic_vector (24 downto 0);	  
	r12 :in std_logic_vector (24 downto 0);
	r13 :in std_logic_vector (24 downto 0);
	r14 :in std_logic_vector (24 downto 0);
	r15 :in std_logic_vector (24 downto 0);
	r16 :in std_logic_vector (24 downto 0);
	r17 :in std_logic_vector (24 downto 0);
	r18 :in std_logic_vector (24 downto 0);
	r19 :in std_logic_vector (24 downto 0);
	r20 :in std_logic_vector (24 downto 0);
	
	r21 :in std_logic_vector (24 downto 0);	  
	r22 :in std_logic_vector (24 downto 0);
	r23 :in std_logic_vector (24 downto 0);
	r24 :in std_logic_vector (24 downto 0);
	r25 :in std_logic_vector (24 downto 0);
	r26 :in std_logic_vector (24 downto 0);
	r27 :in std_logic_vector (24 downto 0);
	r28 :in std_logic_vector (24 downto 0);
	r29 :in std_logic_vector (24 downto 0);
	r30 :in std_logic_vector (24 downto 0);
	
	r31 :in std_logic_vector (24 downto 0);	  
	r32 :in std_logic_vector (24 downto 0);
	r33 :in std_logic_vector (24 downto 0);
	r34 :in std_logic_vector (24 downto 0);
	r35 :in std_logic_vector (24 downto 0);
	r36 :in std_logic_vector (24 downto 0);
	r37 :in std_logic_vector (24 downto 0);
	r38 :in std_logic_vector (24 downto 0);
	r39 :in std_logic_vector (24 downto 0);
	r40 :in std_logic_vector (24 downto 0);		
	
	r41 :in std_logic_vector (24 downto 0);	  
	r42 :in std_logic_vector (24 downto 0);
	r43 :in std_logic_vector (24 downto 0);
	r44 :in std_logic_vector (24 downto 0);
	r45 :in std_logic_vector (24 downto 0);
	r46 :in std_logic_vector (24 downto 0);
	r47 :in std_logic_vector (24 downto 0);
	r48 :in std_logic_vector (24 downto 0);
	r49 :in std_logic_vector (24 downto 0);
	r50 :in std_logic_vector (24 downto 0);
	
	r51 :in std_logic_vector (24 downto 0);	  
	r52 :in std_logic_vector (24 downto 0);
	r53 :in std_logic_vector (24 downto 0);
	r54 :in std_logic_vector (24 downto 0);
	r55 :in std_logic_vector (24 downto 0);
	r56 :in std_logic_vector (24 downto 0);
	r57 :in std_logic_vector (24 downto 0);
	r58 :in std_logic_vector (24 downto 0);
	r59 :in std_logic_vector (24 downto 0);
	r60 :in std_logic_vector (24 downto 0);
	
	r61 :in std_logic_vector (24 downto 0);	  
	r62 :in std_logic_vector (24 downto 0);
	r63 :in std_logic_vector (24 downto 0);
	r64 :in std_logic_vector (24 downto 0);	
	output : out std_logic_vector (24 downto 0)
	);
end instruction_buffer;

--}} End of automatically maintained section

architecture instruction_buffer of instruction_buffer is
type std_logic_aoa is array (0 to 63) of std_logic_vector(24 downto 0);
signal regs : std_logic_aoa;
begin
	
	process(clk)
	begin
		if(rising_edge(clk)) then
			output <= regs(PC);
		end if;
	end process;
	
end instruction_buffer;
